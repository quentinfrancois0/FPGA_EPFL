
module system (
	clk_clk,
	parallel_port0_0_export_0_portp,
	parallel_port0_1_export_0_portp,
	reset_reset_n);	

	input		clk_clk;
	inout	[7:0]	parallel_port0_0_export_0_portp;
	inout	[7:0]	parallel_port0_1_export_0_portp;
	input		reset_reset_n;
endmodule
