
module system (
	clk_clk,
	reset_reset_n,
	pwm_export);	

	input		clk_clk;
	input		reset_reset_n;
	output		pwm_export;
endmodule
